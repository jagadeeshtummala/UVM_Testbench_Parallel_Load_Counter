// package counter_package;
// import uvm_pkg::*;
// `include "uvm_macros.svh"
// `include "packet.sv"
// `include "packet_sequence.sv"
// `include "sequencer.sv"
// `include "driver.sv"
// `include "monitor.sv"
// `include "scoreboard.sv"
// `include "agent.sv"
// `include "environment.sv"

// endpackage : counter_package

`include "uvm_macros.svh"
`include "packet.sv"
`include "packet_sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "environment.sv"